-------------------------------------------------------------------------
-- Joseph Zambreno
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- tb_dff.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a simple VHDL testbench for the
-- edge-triggered flip-flop with parallel access and reset.
--
--
-- NOTES:
-- 8/19/16 by JAZ::Design created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_mux32 is
end tb_mux32;


architecture behavior of tb_mux32 is

component mux32
port(i_1	: in std_logic_vector(31 downto 0);
     i_2	: in std_logic_vector(31 downto 0);
     i_3	: in std_logic_vector(31 downto 0);
     i_4	: in std_logic_vector(31 downto 0);
     i_5	: in std_logic_vector(31 downto 0);
     i_6	: in std_logic_vector(31 downto 0);
     i_7	: in std_logic_vector(31 downto 0);
     i_8	: in std_logic_vector(31 downto 0);
     i_9	: in std_logic_vector(31 downto 0);
     i_10	: in std_logic_vector(31 downto 0);
     i_11	: in std_logic_vector(31 downto 0);
     i_12	: in std_logic_vector(31 downto 0);
     i_13	: in std_logic_vector(31 downto 0);
     i_14	: in std_logic_vector(31 downto 0);
     i_15	: in std_logic_vector(31 downto 0);
     i_16	: in std_logic_vector(31 downto 0);
     i_17	: in std_logic_vector(31 downto 0);
     i_18	: in std_logic_vector(31 downto 0);
     i_19	: in std_logic_vector(31 downto 0);
     i_20	: in std_logic_vector(31 downto 0);
     i_21	: in std_logic_vector(31 downto 0);
     i_22	: in std_logic_vector(31 downto 0);
     i_23	: in std_logic_vector(31 downto 0);
     i_24	: in std_logic_vector(31 downto 0);
     i_25	: in std_logic_vector(31 downto 0);
     i_26	: in std_logic_vector(31 downto 0);
     i_27	: in std_logic_vector(31 downto 0);
     i_28	: in std_logic_vector(31 downto 0);
     i_29	: in std_logic_vector(31 downto 0);
     i_30	: in std_logic_vector(31 downto 0);
     i_31	: in std_logic_vector(31 downto 0);
     i_32	: in std_logic_vector(31 downto 0);
     i_S	: in std_logic_vector(4 downto 0);
     o_F	: out std_logic_vector(31 downto 0));
end component;

signal s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, 
	s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_F	: std_logic_vector(31 downto 0);
signal s_S	: std_logic_vector(4 downto 0);

begin

mux : mux32
port map(i_1 => s_1,
	 i_2 => s_2,
	 i_3 => s_3,
	 i_4 => s_4,
	 i_5 => s_5,
	 i_6 => s_6,
	 i_7 => s_7,
	 i_8 => s_8,
	 i_9 => s_9,
	 i_10 => s_10,
	 i_11 => s_11,
	 i_12 => s_12,
	 i_13 => s_13,
	 i_14 => s_14,
	 i_15 => s_15,
	 i_16 => s_16,
	 i_17 => s_17,
	 i_18 => s_18,
	 i_19 => s_19,
	 i_20 => s_20,
	 i_21 => s_21,
	 i_22 => s_22,
	 i_23 => s_23,
	 i_24 => s_24,
	 i_25 => s_25,
	 i_26 => s_26,
	 i_27 => s_27,
	 i_28 => s_28,
	 i_29 => s_29,
	 i_30 => s_30,
	 i_31 => s_31,
	 i_32 => s_32,
	 o_F => s_F,
	 i_S => s_S);

process
begin

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"00000";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"00001";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"00010";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"00011";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"00100";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"11101";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"11100";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"11011";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"11010";
wait for 100 ns;

s_1 <= x"00000001";
s_2 <= x"00000002";
s_3 <= x"00000004";
s_4 <= x"00000008";
s_5 <= x"00000010";
s_6 <= x"00000020";
s_7 <= x"00000040";
s_8 <= x"00000080";
s_9 <= x"00000100";
s_10 <= x"00000200";
s_11 <= x"00000400";
s_12 <= x"00000800";
s_13 <= x"00001000";
s_14 <= x"00002000";
s_15 <= x"00004000";
s_16 <= x"00008000";
s_17 <= x"00010000";
s_18 <= x"00020000";
s_19 <= x"00040000";
s_20 <= x"00080000";
s_21 <= x"00100000";
s_22 <= x"00200000";
s_23 <= x"00400000";
s_24 <= x"00800000";
s_25 <= x"01000000";
s_26 <= x"02000000";
s_27 <= x"04000000";
s_28 <= x"08000000";
s_29 <= x"10000000";
s_30 <= x"20000000";
s_31 <= x"40000000";
s_32 <= x"80000000";
s_S <= b"11111";
wait for 100 ns;

end process;

end behavior;