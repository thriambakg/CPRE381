    Mac OS X            	   2   �                                           ATTR         �   X                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl   `    �/�8     �; $�J���3Rh�� �Z�ZET�aQ��\��                                    